module FSM_Stop_Watch(
  
);
